// Description: Set global FPGA defines for VCU128
// Author: Vincenzo Maisto vincenzo.maisto2@unina.it

`define xcvu37p
